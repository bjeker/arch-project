module not_4b(x, out);

  output [3:0] out, o;
  input [3:0] x;

  wire x, out;

  assign out = ~x;

endmodule