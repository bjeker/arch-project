module shift_4b(x, y);

  output xOut, yOut;
  input x, y;

  wire x, y, xOut, yOut;

  assign xOut = x;
  assign yOut = y;

endmodule