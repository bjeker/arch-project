module xor_4b(x, y, out);

  output [3:0] out;
  input [3:0] x, y;

  wire x, y, out;

  assign out = x ^ y;

endmodule
