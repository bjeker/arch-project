module shift_4b(x, y);

  output [3:0] xOut, yOut;
  input [3:0] x, y;

  wire [3:0] x, y, xOut, yOut;

  assign xOut = x;
  assign yOut = y;

endmodule