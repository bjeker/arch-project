module shift_4b(x);

  output out;
  input x;

  wire x, out;

  assign out = x;

endmodule
