module not_1b(x, out);

  output out;
  input x;

  wire x, out;

  assign out = ~x;

endmodule
